module top_module(
    input a,
    input b,
    input c,
    output out  ); 

    or(out, a, b, c);
endmodule
